module mce(a, b, max, min);
    input logic [7:0] a;
    input logic [7:0] b;

    output logic [7:0] max;
    output logic [7:0] min;

endmodule:mce
