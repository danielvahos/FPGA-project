module vga(
    input wire pixel_clk,
    input wire pixel_rst,
    video_if.master video_ifm
);
